package l1_cache_types;

typedef logic [127:0] l1_cache_line
typedef logic [9:0]   l1_cache_tag       

endpackage : l1_cache_types
