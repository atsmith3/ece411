package lc3b_ctypes;

typedef logic [127:0] lc3b_cline;
typedef logic [8:0]   lc3b_ctag;
typedef logic [2:0]   lc3b_cindex;
typedef logic [3:0]   lc3b_coffset;

endpackage : lc3b_ctypes
