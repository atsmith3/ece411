import ../lc3b_types::*;
import lc3b_cache_types::*;

module cache
(
   input logic clk,

   /* Input Logic (from LC3) */
   lc3b_word 
);



endmodule : cache
